--
-- Notes on using `gtu-pkgpatch-ipbus' for this package:
--  * _IPBUS_TIMESTAMP_    32 bit UNIX timestamp placeholder (X"00000000")
--  * _IPBUS_USERNAME_     unix username 32 char string placeholder (X"...")
--  * _IPBUS_HOSTNAME_     machine hostname 32 char string placeholder (X"...")
--
--------------------------------------------------------------------------------

library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.top_decl.all;

package gt_top_pkg is

-- BA 2014-08-06: TIMESTAMP generated by gtu-pkgpatch-ipbus (32 bits), has to be interpreted as 32 bit UNIX timestamp.
constant TOP_TIMESTAMP : std_logic_vector(31 downto 0) := X"59A81F11";
-- HB 2014-05-23: USERNAME generated by gtu-pkgpatch-ipbus (256 bits = 8 x 32 bits), has to be interpreted as 32 ASCII-characters string (from right to left).
constant TOP_USERNAME : std_logic_vector(32*8-1 downto 0)  := X"0000000000000000000000000000000000000000000000007265756167726562";
-- HB 2014-05-23: HOSTNAME generated by gtu-pkgpatch-ipbus (256 bits = 8 x 32 bits), has to be interpreted as 32 ASCII-characters string (from right to left).
constant TOP_HOSTNAME : std_logic_vector(32*8-1 downto 0) := X"00000000000000000000000000000000000000000000000000326163746d7467";

end;



