-- Description:
-- Global Trigger Logic module.

-- HB 2019-06-27: Changed type of conversion signals.
-- HB 2019-03-08: new strcture with instance of l1menu.vhd

library ieee;
use ieee.std_logic_1164.all;

use work.gtl_pkg.all;
use work.l1menu_pkg.ALL;

entity gtl_module is
    port(
        lhc_clk : in std_logic;
        data_in : in gtl_data_record;
        algo_o : out std_logic_vector(NR_ALGOS-1 downto 0));
end gtl_module;

architecture rtl of gtl_module is
    
    signal data_p : data_pipeline_record;
    signal conv : conv_pipeline_record;
    signal algo : std_logic_vector(NR_ALGOS-1 downto 0) := (others => '0');

begin

-- +/-2 BX pipeline for input data and conversions of object parameters
    bx_pipeline_i: entity work.bx_pipeline
        port map(
            lhc_clk, data_in, data_p, conv
        );

-- Module l1menu.vhd contains VHDL representation of L1Menu,
-- generated by VHDL Producer
    l1menu_i: entity work.l1menu
        port map(
            lhc_clk, data_p, conv, algo
        );

-- Pipeline stages for algorithms
    algo_pipeline_i: entity work.delay_pipeline
        generic map(
            DATA_WIDTH => NR_ALGOS,
            STAGES => ALGO_REG_STAGES
        )
        port map(
            lhc_clk, algo, algo_o
        );

end architecture rtl;
